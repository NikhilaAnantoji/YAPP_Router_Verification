package yapp_pkg;

  // import the UVM library
  import uvm_pkg::*;

  // include the UVM macros
  `include "uvm_macros.svh"

  // include the YAPP packet definition
  `include "yapp.svh"

endpackage : yapp_pkg
